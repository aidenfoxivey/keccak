library ieee;
use ieee.std_logic_1164.all;

library work;
use work.keccak_common.all;

-- https://keccak.team/keccak_specs_summary.html
package keccak_constants is
    type round_constant_array_t is array (0 to 23) of lane;

    constant ROUND_CONSTANTS : round_constant_array_t
     := (
        0 => X"0000000000000001",
        1 => X"0000000000008082",
        2 => X"800000000000808A",
        3 => X"8000000080008000",
        4 => X"000000000000808B",
        5 => X"0000000080000001",
        6 => X"8000000080008081",
        7 => X"8000000000008009",
        8 => X"000000000000008A",
        9 => X"0000000000000088",
        10 => X"0000000080008009",
        11 => X"000000008000000A",
        12 => X"000000008000808B",
        13 => X"800000000000008B",
        14 => X"8000000000008089",
        15 => X"8000000000008003",
        16 => X"8000000000008002",
        17 => X"8000000000000080",
        18 => X"000000000000800A",
        19 => X"800000008000000A",
        20 => X"8000000080008081",
        21 => X"8000000000008080",
        22 => X"0000000080000001",
        23 => X"8000000080008008"
    );

    type rotation_offsets_t is array (0 to 4, 0 to 4) of natural;

    constant ROTATION_OFFSETS : rotation_offsets_t := (
        -- x = 0 (y = 0,1,2,3,4)
        (0 => 0, 1 => 36, 2 => 3, 3 => 41, 4 => 18),
        -- x = 1 (y = 0,1,2,3,4)
        (0 => 1, 1 => 44, 2 => 10, 3 => 45, 4 => 2),
        -- x = 2 (y = 0,1,2,3,4)
        (0 => 62, 1 => 6, 2 => 43, 3 => 15, 4 => 61),
        -- x = 3 (y = 0,1,2,3,4)
        (0 => 28, 1 => 55, 2 => 25, 3 => 21, 4 => 56),
        -- x = 4 (y = 0,1,2,3,4)
        (0 => 27, 1 => 20, 2 => 39, 3 => 8, 4 => 14)
    );

end package keccak_constants;
